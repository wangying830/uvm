module m2;
  initial begin
    $display("This is dummy m2");
  end
endmodule
