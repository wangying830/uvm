module m1;
  m2 m2_inst();
endmodule
