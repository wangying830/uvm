module top;
  m1 m1_inst();
endmodule
