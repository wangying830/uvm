// timescale = 1ps/1ps
// default delay
int PORT0_DELAY = 1000;
int PORT1_DELAY = 1100;
int PORT2_DELAY = 1200;
int PORT3_DELAY = 1300;
int PORT4_DELAY = 1400;

