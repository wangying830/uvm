module m2;
  logic v1, v2;
  initial begin
    $display("This is m2");
  end
endmodule
